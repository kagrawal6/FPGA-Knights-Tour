//`timescale 1ns/1ps
module Knights_Post_Synth_tb();
	import  tb_tasks::*;

	localparam FAST_SIM = 1;


	/////////////////////////////
	// Stimulus of type reg //
	/////////////////////////
	reg clk, RST_n;
	reg [15:0] cmd;
	reg send_cmd;

	///////////////////////////////////
	// Declare any internal signals //
	/////////////////////////////////
	wire SS_n,SCLK,MOSI,MISO,INT;
	wire lftPWM1,lftPWM2,rghtPWM1,rghtPWM2;
	wire TX_RX, RX_TX;
	logic cmd_sent;
	logic resp_rdy;
	logic [7:0] resp;
	wire IR_en;
	wire lftIR_n,rghtIR_n,cntrIR_n;

	//////////////////////
	// Instantiate DUT //
	////////////////////
	KnightsTour iDUT(.clk(clk), .RST_n(RST_n), .SS_n(SS_n), .SCLK(SCLK),
					.MOSI(MOSI), .MISO(MISO), .INT(INT), .lftPWM1(lftPWM1),
					.lftPWM2(lftPWM2), .rghtPWM1(rghtPWM1), .rghtPWM2(rghtPWM2),
					.RX(TX_RX), .TX(RX_TX), .piezo(piezo), .piezo_n(piezo_n),
					.IR_en(IR_en), .lftIR_n(lftIR_n), .rghtIR_n(rghtIR_n),
					.cntrIR_n(cntrIR_n));
					
	/////////////////////////////////////////////////////
	// Instantiate RemoteComm to send commands to DUT //
	///////////////////////////////////////////////////
	RemoteComm iRMT(.clk(clk), .rst_n(RST_n), .RX(RX_TX), .TX(TX_RX), .cmd(cmd),
				.snd_cmd(send_cmd), .cmd_snt(cmd_sent), .resp_rdy(resp_rdy), .resp(resp));
					
	//////////////////////////////////////////////////////
	// Instantiate model of Knight Physics (and board) //
	////////////////////////////////////////////////////
	KnightPhysics iPHYS(.clk(clk),.RST_n(RST_n),.SS_n(SS_n),.SCLK(SCLK),.MISO(MISO),
						.MOSI(MOSI),.INT(INT),.lftPWM1(lftPWM1),.lftPWM2(lftPWM2),
						.rghtPWM1(rghtPWM1),.rghtPWM2(rghtPWM2),.IR_en(IR_en),
						.lftIR_n(lftIR_n),.rghtIR_n(rghtIR_n),.cntrIR_n(cntrIR_n)); 

    initial begin
        clk = 0;
        RST_n = 0;
        
        send_cmd = 0;
        
        @(negedge clk);
        RST_n = 1;
        repeat(1000000)@(posedge clk);
        @(negedge clk);
        cmd = 15'h2000;
        
        // Pulsing send_cmd
        @(negedge clk);
        send_cmd = 1;
        
        @(negedge clk);
        send_cmd = 0;

        repeat(1000000)@(posedge clk);
        SendCmd(.host_cmd(16'h4002),.cmd(cmd), .send_cmd(send_cmd),.clk(clk));
        @(posedge resp_rdy);
        repeat(1000000)@(posedge clk);
        $stop();
    end
    always  
        #5 clk= ~clk;
endmodule